    `include "axis_data.svh"
    
    `include "axis_sequence_config.svh"
    `include "axis_sequence.svh"
    
    `include "axis_sequencer.svh"
    `include "axis_driver.svh"
    `include "axis_monitor.svh"

    `include "axis_agent.svh"
