package test_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "../../src/axis_include.svh"

    `include "test_env.svh"
    `include "rand_axis_test.svh"
    
endpackage